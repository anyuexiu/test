module AXI_waddr(
	aclk,
	areset,
	//
);

input aclk;
input areset;


endmodule
